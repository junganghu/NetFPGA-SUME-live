//
// Copyright (C) 2015 Digilent Inc.
// All rights reserved.
//
// @NETFPGA_LICENSE_HEADER_START@
//
// Licensed to NetFPGA C.I.C. (NetFPGA) under one or more contributor
// license agreements.  See the NOTICE file distributed with this work for
// additional information regarding copyright ownership.  NetFPGA licenses this
// file to you under the NetFPGA Hardware-Software License, Version 1.0 (the
// "License"); you may not use this file except in compliance with the
// License.  You may obtain a copy of the License at:
//
//   http://www.netfpga-cic.org
//
// Unless required by applicable law or agreed to in writing, Work distributed
// under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
//
// @NETFPGA_LICENSE_HEADER_END@
//

`timescale 1 ps / 1 ps

	module nf_sume_gpio_test #
	(
		// Users to add parameters here

		// User parameters ends
		// Do not modify the parameters beyond this line


		// Parameters of Axi Slave Bus Interface S_AXI
		parameter integer C_S_AXI_DATA_WIDTH	= 32,
		parameter integer C_S_AXI_ADDR_WIDTH	= 5
	)
	(
		// Users to add ports here
		inout wire [33:0] fmc_la_odd,
		inout wire [33:0] fmc_la_even,
		inout wire [3:0] pmod_up,
		inout wire [3:0] pmod_down,
		output wire [3:0] pmod_up_dir,
		output wire [3:0] pmod_down_dir,
		output wire pmod_oe,
		// User ports ends
		// Do not modify the ports beyond this line

		// Ports of Axi Slave Bus Interface S_AXI
		input wire  s_axi_aclk,
		input wire  s_axi_aresetn,
		input wire [C_S_AXI_ADDR_WIDTH-1 : 0] s_axi_awaddr,
		input wire [2 : 0] s_axi_awprot,
		input wire  s_axi_awvalid,
		output wire  s_axi_awready,
		input wire [C_S_AXI_DATA_WIDTH-1 : 0] s_axi_wdata,
		input wire [(C_S_AXI_DATA_WIDTH/8)-1 : 0] s_axi_wstrb,
		input wire  s_axi_wvalid,
		output wire  s_axi_wready,
		output wire [1 : 0] s_axi_bresp,
		output wire  s_axi_bvalid,
		input wire  s_axi_bready,
		input wire [C_S_AXI_ADDR_WIDTH-1 : 0] s_axi_araddr,
		input wire [2 : 0] s_axi_arprot,
		input wire  s_axi_arvalid,
		output wire  s_axi_arready,
		output wire [C_S_AXI_DATA_WIDTH-1 : 0] s_axi_rdata,
		output wire [1 : 0] s_axi_rresp,
		output wire  s_axi_rvalid,
		input wire  s_axi_rready
	);
	
    wire [33:0] fmc_gpio_out;
    wire [33:0] fmc_gpio_in;
    wire [3:0] pmod_gpio_out;
    wire [3:0] pmod_gpio_in;
    wire tri_ctrl;
		
// Instantiation of Axi Bus Interface S_AXI
	nf_sume_gpio_test_S_AXI # ( 
		.C_S_AXI_DATA_WIDTH(C_S_AXI_DATA_WIDTH),
		.C_S_AXI_ADDR_WIDTH(C_S_AXI_ADDR_WIDTH)
	) nf_sume_gpio_test_S_AXI_inst (
	    .fmc_gpio_out(fmc_gpio_out),
	    .fmc_gpio_in(fmc_gpio_in),
	    .pmod_gpio_out(pmod_gpio_out),
	    .pmod_gpio_in(pmod_gpio_in),
	    .tri_ctrl(tri_ctrl),
		.S_AXI_ACLK(s_axi_aclk),
		.S_AXI_ARESETN(s_axi_aresetn),
		.S_AXI_AWADDR(s_axi_awaddr),
		.S_AXI_AWPROT(s_axi_awprot),
		.S_AXI_AWVALID(s_axi_awvalid),
		.S_AXI_AWREADY(s_axi_awready),
		.S_AXI_WDATA(s_axi_wdata),
		.S_AXI_WSTRB(s_axi_wstrb),
		.S_AXI_WVALID(s_axi_wvalid),
		.S_AXI_WREADY(s_axi_wready),
		.S_AXI_BRESP(s_axi_bresp),
		.S_AXI_BVALID(s_axi_bvalid),
		.S_AXI_BREADY(s_axi_bready),
		.S_AXI_ARADDR(s_axi_araddr),
		.S_AXI_ARPROT(s_axi_arprot),
		.S_AXI_ARVALID(s_axi_arvalid),
		.S_AXI_ARREADY(s_axi_arready),
		.S_AXI_RDATA(s_axi_rdata),
		.S_AXI_RRESP(s_axi_rresp),
		.S_AXI_RVALID(s_axi_rvalid),
		.S_AXI_RREADY(s_axi_rready)
	);

	// Add user logic here
    // tri_ctrl = 1: FMC_LA_Even - output; FMC_LA_Odd - Input; Pmod_Down - output; Pmod_Up - input
    assign fmc_la_even = (tri_ctrl == 1'b1) ? fmc_gpio_out : 'bz;
    assign fmc_la_odd = (tri_ctrl == 1'b0) ? fmc_gpio_out : 'bz;
    
    assign pmod_down = (tri_ctrl == 1'b1) ? pmod_gpio_out : 'bz;
    assign pmod_up = (tri_ctrl == 1'b0) ? pmod_gpio_out : 'bz;
    
    assign fmc_gpio_in = (tri_ctrl == 1'b1) ? fmc_la_odd : fmc_la_even;
    assign pmod_gpio_in = (tri_ctrl == 1'b1) ? pmod_up : pmod_down;
    
    assign pmod_down_dir = {tri_ctrl, tri_ctrl, tri_ctrl, tri_ctrl};
    assign pmod_up_dir = {~tri_ctrl, ~tri_ctrl, ~tri_ctrl, ~tri_ctrl}; 
    
    assign pmod_oe = 1'b0;
	// User logic ends

	endmodule
